module NOT_Gate (
  input X,
  output Z
);
  assign Z = ~ X;
endmodule 