module Or_Gate (
  input A,
  input B,
  output O
);
  assign O = A|B;

endmodule 