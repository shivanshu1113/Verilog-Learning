module XOR_Gate (
    input A,
    input B,
    output C
);
    assign C = A ^ B;
endmodule